`include"uvm_pkg.sv"
import uvm_pkg::*;
`include"axi_interface.sv"
`include"axi_tx.sv"
`include"axi_sequence.sv"
`include"axi_sequencer.sv"
`include"axi_master_driver.sv"
`include"axi_monitor.sv"
`include"axi_coverage.sv"
`include"axi_scoreboard.sv"
`include"axi_master_agent.sv"
`include"axi_slave_driver.sv"
`include"axi_slave_agent.sv"
`include"axi_master_env.sv"
`include"axi_slave_env.sv"
`include"axi_top_env.sv"
`include"axi_test.sv"
`include"axi_top.sv"
