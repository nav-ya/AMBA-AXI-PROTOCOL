interface axi_interface(input bit aclk,aresetn);
	 logic[7:0] awid;
	 logic awvalid;
	 logic[3:0] awlen;
         logic awready;
	 logic[3:0]awcache;
	 logic[3:0]awsize;
	 logic[1:0]awburst;
	 logic[1:0]awlock;
	 logic[3:0]awprot;
         logic wvalid;
	 logic wready;
         logic[7:0]wid;
         logic[31:0] wdata;
         logic[3:0] wstrb;        
	 logic wlast;
         logic bvalid;
	 logic bready;
         logic[7:0]bid;
         logic[1:0] bresp;
	 logic[31:0] araddr;
	 logic[7:0] arid;
	 logic arvalid;
	 logic[3:0] arlen;
         logic  arready;
	 logic[3:0]arcache;
	 logic[3:0]arsize;
	 logic[1:0]arburst;
	 logic[1:0]arlock;
	 logic[3:0]arprot;         
	 logic rvalid;
	 logic rready;
         logic[7:0]rid;
         logic[31:0] rdata;
	 logic rlast;
	 logic[1:0] rresp;
 endinterface
